module INST_MEM (
    input [63:0] PC,
    input reset,
    output [63:0] command_code
);

    reg [7:0] 
    
endmodule: